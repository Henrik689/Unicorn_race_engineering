-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Tuesday, June 30, 2009 19:05:45 Rom, sommertid

